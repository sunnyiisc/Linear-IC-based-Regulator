*
.tran 50us 100ms uic
.include ic_regulator.net
